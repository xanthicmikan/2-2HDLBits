module top_module( 
    input [255:0] in,
    input [7:0] sel,
    output out );
    
	// Select one bit from vector in[]. The bit being selected can be variable.
    assign out = in[sel]; 

endmodule